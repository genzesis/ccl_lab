** Profile: "SCHEMATIC1-sim2"  [ D:\krishnendu147\rlc-SCHEMATIC1-sim2.sim ] 

** Creating circuit file "rlc-SCHEMATIC1-sim2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 0.5u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rlc-SCHEMATIC1.net" 


.END
