** Profile: "SCHEMATIC1-rlc"  [ D:\krishnendu147\rlc-SCHEMATIC1-rlc.sim ] 

** Creating circuit file "rlc-SCHEMATIC1-rlc.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rlc-SCHEMATIC1.net" 


.END
