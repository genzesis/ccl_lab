** Profile: "SCHEMATIC1-introsim"  [ D:\krishnendu147\introduction-SCHEMATIC1-introsim.sim ] 

** Creating circuit file "introduction-SCHEMATIC1-introsim.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 2ms 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\introduction-SCHEMATIC1.net" 


.END
